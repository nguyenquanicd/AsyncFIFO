//================================================================================
// File name:   asyn_fifo_parameters.vh
// Project:     LAB 5:  Asynchronous FIFO
//Author:   
//================================================================================

    parameter   DATA_WIDTH = 8;
    parameter   POINTER_WIDTH = 3;
    parameter    FIFO_DEPTH = 2**POINTER_WIDTH;
    