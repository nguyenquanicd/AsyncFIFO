//=========================================================================
// File name:   asyn_fifo_define.vh
// Project:     LAB 5: Asynchronous FIFO
// Author:  
//=========================================================================

`define     EMPTY_FLAG;
`define     FULL_FLAG;
`define     OVERFLOW_FLAG;
`define     UNDERFLOW_FLAG;